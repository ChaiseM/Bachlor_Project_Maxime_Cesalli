--
-- VHDL Architecture Splitter.HighLevel.HighLevel
--
-- Created:
--          by - maxime.cesalli.UNKNOWN (WE2330804)
--          at - 14:12:04 14.07.2023
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE HighLevel OF HighLevel IS
BEGIN
    writeEnA <= '1'; 
    writeENB <= '0';
    dataInB <= "0000000000000000";
END ARCHITECTURE HighLevel;

